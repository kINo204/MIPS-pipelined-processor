// alu.vh

localparam  SLL = 4'b0000,
            SRL = 4'b0001,
            SRA = 4'b0010,
            ADD = 4'b0011,
            SUB = 4'b0100,
            AND = 4'b0101,
            OR  = 4'b0110;
// ExcCode
localparam
    EXC_INT  = 0,
    EXC_ADEL = 4,
    EXC_ADES = 5,
    EXC_SYSC = 8,
    EXC_RIST = 10,
    EXC_OVFL = 12;
// mudv.vh

localparam  TIME_MUL = 5,
            TIME_DIV = 10;

localparam  MULT  = 3'b000,
            MULTU = 3'b001,
            DIV   = 3'b010,
            DIVU  = 3'b011,
            MDSP  = 3'b100;